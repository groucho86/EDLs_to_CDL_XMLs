<?xml version="1.0" ?>
<ColorDecisionList>
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Slope>1.376302 1.350373 1.156858</Slope>
				<Offset>-0.061675 -0.074797 -0.024712</Offset>
				<Power>1.532946 1.548055 1.533721</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.000000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
