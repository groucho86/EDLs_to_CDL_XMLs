<?xml version="1.0" ?>
<ColorDecisionList>
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Slope>1.796064 1.554420 1.498708</Slope>
				<Offset>-0.161735 -0.044558 0.058580</Offset>
				<Power>2.098053 1.959595 2.020724</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.000000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
