<?xml version="1.0" ?>
<ColorDecisionList>
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Slope>1.153253 1.091636 1.106670</Slope>
				<Offset>0.146810 0.138966 0.140880</Offset>
				<Power>3.241508 3.256578 3.255717</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.000000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
