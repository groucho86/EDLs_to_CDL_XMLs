<?xml version="1.0" ?>
<ColorDecisionList>
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Slope>1.887539 1.896713 1.869297</Slope>
				<Offset>-0.146187 -0.143821 -0.175531</Offset>
				<Power>1.355141 1.279595 1.475515</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.000000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
