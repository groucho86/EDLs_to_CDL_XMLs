<?xml version="1.0" ?>
<ColorDecisionList>
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Slope>1.286208 1.203307 1.217375</Slope>
				<Offset>0.147690 0.210024 0.164590</Offset>
				<Power>3.964272 3.615482 3.934752</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.000000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
