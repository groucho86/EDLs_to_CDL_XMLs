<?xml version="1.0" ?>
<ColorDecisionList>
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Slope>1.876222 1.545198 1.286441</Slope>
				<Offset>-0.431919 -0.225799 -0.012615</Offset>
				<Power>2.502286 2.504979 2.493689</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.000000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
