<?xml version="1.0" ?>
<ColorDecisionList>
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Slope>1.564273 1.324745 1.287985</Slope>
				<Offset>-0.143760 -0.007883 0.060659</Offset>
				<Power>2.266541 2.264585 2.255546</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.000000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
