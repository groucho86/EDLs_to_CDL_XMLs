<?xml version="1.0" ?>
<ColorDecisionList>
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Slope>1.752198 1.563238 1.099331</Slope>
				<Offset>-0.205091 -0.070173 -0.112716</Offset>
				<Power>1.910205 1.910205 1.910205</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.000000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
