<?xml version="1.0" ?>
<ColorDecisionList>
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Slope>1.859397 1.721146 1.590698</Slope>
				<Offset>-0.180457 -0.167040 -0.154380</Offset>
				<Power>1.703328 1.703328 1.703551</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.000000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
