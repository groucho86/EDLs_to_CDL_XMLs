<?xml version="1.0" ?>
<ColorDecisionList>
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Slope>1.110770 1.079979 1.169953</Slope>
				<Offset>0.032561 0.019570 -0.011226</Offset>
				<Power>1.841824 1.910732 1.913079</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.000000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
