<?xml version="1.0" ?>
<ColorDecisionList>
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Slope>1.197091 1.178911 1.276364</Slope>
				<Offset>0.018709 0.005404 -0.029054</Offset>
				<Power>1.898249 1.969163 1.971382</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.000000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
